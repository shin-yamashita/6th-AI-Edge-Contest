
package pkg_rv_decode;

`include "rv_exp_cinsn.sv"      // C-insn expand table
`include "rv_dec_insn.sv"       // insn decode table 

endpackage


