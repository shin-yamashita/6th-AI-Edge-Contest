//
// logic type deffs
//

`ifndef RV_TYPES_H
`define RV_TYPES_H

 typedef logic [1:0]         u2_t;
 typedef logic [2:0]         u3_t;
 typedef logic [3:0]         u4_t;
 typedef logic [4:0]         u5_t;
 typedef logic [5:0]         u6_t;
 typedef logic [6:0]         u7_t;
 typedef logic [7:0]         u8_t;
 typedef logic signed [7:0]  s8_t;
 typedef logic [8:0]         u9_t;
 typedef logic [11:0]        u12_t;
 typedef logic signed [11:0] s12_t;
 typedef logic [15:0]        u16_t;
 typedef logic signed [15:0] s16_t;
 typedef logic [16:0]        u17_t;
 typedef logic signed [16:0] s17_t;
 typedef logic [19:0]        u20_t;
 typedef logic [21:0]        u22_t;
 typedef logic [23:0]        u24_t;
 typedef logic signed [23:0] s24_t;
 typedef logic [25:0]        u26_t;
 typedef logic [26:0]        u27_t;
 typedef logic [27:0]        u28_t;
 typedef logic [28:0]        u29_t;
 typedef logic [31:0]        u32_t;
 typedef logic signed [31:0] s32_t;
 typedef logic [32:0]        u33_t;
 typedef logic signed [32:0] s33_t;
 typedef logic [33:0]        u34_t;
 typedef logic signed [33:0] s34_t;
 typedef logic [47:0]        u48_t;
 typedef logic [63:0]        u64_t;
 typedef logic signed [63:0] s64_t;

`endif

